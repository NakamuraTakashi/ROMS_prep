netcdf Yaeyama1_river_v3 {
dimensions:
	xi_rho = 310 ;
	xi_u = 309 ;
	xi_v = 310 ;
	eta_rho = 280 ;
	eta_u = 280 ;
	eta_v = 279 ;
	s_rho = 30 ;
	river = 5 ;
	river_time = 20 ;
variables:
	double river(river) ;
		river:long_name = "river runoff identification number" ;
	double river_Xposition(river) ;
		river_Xposition:long_name = "river XI-position at RHO-points" ;
		river_Xposition:valid_min = 1. ;
		river_Xposition:valid_max = 309. ;
	double river_Eposition(river) ;
		river_Eposition:long_name = "river ETA-position at RHO-points" ;
		river_Eposition:valid_min = 1. ;
		river_Eposition:valid_max = 279. ;
	double river_direction(river) ;
		river_direction:long_name = "river runoff direction" ;
	double river_Vshape(s_rho, river) ;
		river_Vshape:long_name = "river runoff mass transport vertical profile" ;
	double river_time(river_time) ;
		river_time:long_name = "river runoff time" ;
		river_time:units = "days since 2014-04-01 00:00:00" ;
		river_time:add_offset = 0. ;
	double river_transport(river_time, river) ;
		river_transport:long_name = "river runoff vertically integrated mass transport" ;
		river_transport:units = "meter3 second-1" ;
		river_transport:time = "river_time" ;
	double river_temp(river_time, s_rho, river) ;
		river_temp:long_name = "river runoff potential temperature" ;
		river_temp:units = "Celsius" ;
		river_temp:time = "river_time" ;
	double river_salt(river_time, s_rho, river) ;
		river_salt:long_name = "river runoff salinity" ;
		river_salt:time = "river_time" ;

// global attributes:
		:type = "ROMS FORCING file" ;
		:title = "YAEYAMA River Forcing" ;
		:grd_file = "Yaeyama1_grd_v8.nc" ;
		:rivers = "(1)Nakama river, (2) Nagra river, (3) Arakawa river, (4) Miyara river, (5) Todoroki river" ;
data:

 river = 1, 2, 3, 4, 5 ;

 river_Xposition = 74, 191, 191, 196, 199 ;

 river_Eposition = 82, 91, 87, 89, 91 ;

 river_direction = 0, 0, 0, 1, 0 ;

 river_Vshape =
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0.005, 0.005, 0.005, 0.005, 0.005,
  0.005, 0.005, 0.005, 0.005, 0.005,
  0.005, 0.005, 0.005, 0.005, 0.005,
  0.005, 0.005, 0.005, 0.005, 0.005,
  0.005, 0.005, 0.005, 0.005, 0.005,
  0.005, 0.005, 0.005, 0.005, 0.005,
  0.01, 0.01, 0.01, 0.01, 0.01,
  0.01, 0.01, 0.01, 0.01, 0.01,
  0.01, 0.01, 0.01, 0.01, 0.01,
  0.01, 0.01, 0.01, 0.01, 0.01,
  0.02, 0.02, 0.02, 0.02, 0.02,
  0.02, 0.02, 0.02, 0.02, 0.02,
  0.02, 0.02, 0.02, 0.02, 0.02,
  0.02, 0.02, 0.02, 0.02, 0.02,
  0.03, 0.03, 0.03, 0.03, 0.03,
  0.03, 0.03, 0.03, 0.03, 0.03,
  0.03, 0.03, 0.03, 0.03, 0.03,
  0.04, 0.04, 0.04, 0.04, 0.04,
  0.04, 0.04, 0.04, 0.04, 0.04,
  0.04, 0.04, 0.04, 0.04, 0.04,
  0.05, 0.05, 0.05, 0.05, 0.05,
  0.06, 0.06, 0.06, 0.06, 0.06,
  0.07, 0.07, 0.07, 0.07, 0.07,
  0.08, 0.08, 0.08, 0.08, 0.08,
  0.09, 0.09, 0.09, 0.09, 0.09,
  0.09, 0.09, 0.09, 0.09, 0.09,
  0.1, 0.1, 0.1, 0.1, 0.1,
  0.1, 0.1, 0.1, 0.1, 0.1 ;

 river_time = 0, 15, 30, 45, 60, 75, 90, 105, 120, 135, 150, 165, 180, 195, 
    210, 225, 240, 255, 270, 285 ;

 river_transport =
  50, -20, -5, -20, 1,
  50, -20, -5, -20, 1,
  50, -20, -5, -20, 1,
  50, -20, -5, -20, 1,
  50, -20, -5, -20, 1,
  50, -20, -5, -20, 1,
  50, -20, -5, -20, 1,
  50, -20, -5, -20, 1,
  50, -20, -5, -20, 1,
  50, -20, -5, -20, 1,
  50, -20, -5, -20, 1,
  50, -20, -5, -20, 1,
  50, -20, -5, -20, 1,
  50, -20, -5, -20, 1,
  50, -20, -5, -20, 1,
  50, -20, -5, -20, 1,
  50, -20, -5, -20, 1,
  50, -20, -5, -20, 1,
  50, -20, -5, -20, 1,
  50, -20, -5, -20, 1 ;

 river_temp =
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20,
  20, 20, 20, 20, 20 ;

 river_salt =
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0 ;
}
