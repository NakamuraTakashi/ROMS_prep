netcdf TokyoBay3_river_2d_2018_2020 {
dimensions:
    s_rho = 30 ;
	river = 9 ;
	river_time = UNLIMITED ; // (0 currently)
variables:
	double river(river) ;
		river:long_name = "river runoff identification number" ;
	double river_Xposition(river) ;
		river_Xposition:long_name = "river XI-position" ;
		river_Xposition:LuvSrc_meaning = "i point index of U or V face source/sink" ;
		river_Xposition:LwSrc_meaning = "i point index of RHO center source/sink" ;
	double river_Eposition(river) ;
		river_Eposition:long_name = "river ETA-position" ;
		river_Eposition:LuvSrc_meaning = "j point index of U or V face source/sink" ;
		river_Eposition:LwSrc_meaning = "j point index of RHO center source/sink" ;
	double river_direction(river) ;
		river_direction:long_name = "river runoff direction" ;
		river_direction:flag_values = "0, 1" ;
		river_direction:flag_meanings = "flow across u-face, flow across v-face" ;
		river_direction:LwSrc_True = "flag not used" ;
	double river_Vshape(s_rho, river) ;
		river_Vshape:long_name = "river runoff mass transport vertical profile" ;
		river_Vshape:requires = "must sum to 1 over s_rho" ;
	double river_time(river_time) ;
		river_time:long_name = "river runoff time" ;
		river_time:units = "days since 2000-01-01 00:00:00" ;
	double river_transport(river_time, river) ;
		river_transport:long_name = "river runoff vertically integrated mass transport" ;
		river_transport:units = "meter3 second-1" ;
		river_transport:time = "river_time" ;
	double river_salt(river_time, river) ;
		river_salt:long_name = "river runoff salinity" ;
		river_salt:time = "river_time" ;
	double river_temp(river_time, river) ;
		river_temp:long_name = "river runoff potential temperature" ;
		river_temp:units = "Celsius" ;
		river_temp:time = "river_time" ;
	double river_DO(river_time, river) ;
		river_DO:long_name = "river runoff DO" ;
		river_DO:units = "umol L-1" ;
		river_DO:time = "river_time" ;
	double river_TA(river_time, river) ;
		river_TA:long_name = "river runoff alkalinity" ;
		river_TA:units = "umol kg-1" ;
		river_TA:time = "river_time" ;
	double river_DIC_01(river_time, river) ;
		river_DIC_01:long_name = "river runoff DIC_01" ;
		river_DIC_01:units = "umol kg-1" ;
		river_DIC_01:time = "river_time" ;
	double river_NO3_01(river_time, river) ;
		river_NO3_01:long_name = "river runoff NO3_01" ;
		river_NO3_01:units = "umol L-1" ;
		river_NO3_01:time = "river_time" ;
	double river_NH4_01(river_time, river) ;
		river_NH4_01:long_name = "river runoff NH4_01" ;
		river_NH4_01:units = "umol L-1" ;
		river_NH4_01:time = "river_time" ;
	double river_PO4_01(river_time, river) ;
		river_PO4_01:long_name = "river runoff PO4_01" ;
		river_PO4_01:units = "umol L-1" ;
		river_PO4_01:time = "river_time" ;
	double river_DOC01_01(river_time, river) ;
		river_DOC01_01:long_name = "river runoff DOC01_01" ;
		river_DOC01_01:units = "umol L-1" ;
		river_DOC01_01:time = "river_time" ;
	double river_DOC02_01(river_time, river) ;
		river_DOC02_01:long_name = "river runoff DOC02_01" ;
		river_DOC02_01:units = "umol L-1" ;
		river_DOC02_01:time = "river_time" ;
	double river_DON01_01(river_time, river) ;
		river_DON01_01:long_name = "river runoff DON01_01" ;
		river_DON01_01:units = "umol L-1" ;
		river_DON01_01:time = "river_time" ;
	double river_DON02_01(river_time, river) ;
		river_DON02_01:long_name = "river runoff DON02_01" ;
		river_DON02_01:units = "umol L-1" ;
		river_DON02_01:time = "river_time" ;
	double river_DOP01_01(river_time, river) ;
		river_DOP01_01:long_name = "river runoff DOP01_01" ;
		river_DOP01_01:units = "umol L-1" ;
		river_DOP01_01:time = "river_time" ;
	double river_DOP02_01(river_time, river) ;
		river_DOP02_01:long_name = "river runoff DOP02_01" ;
		river_DOP02_01:units = "umol L-1" ;
		river_DOP02_01:time = "river_time" ;
	double river_POC01_01(river_time, river) ;
		river_POC01_01:long_name = "river runoff POC01_01" ;
		river_POC01_01:units = "umol L-1" ;
		river_POC01_01:time = "river_time" ;
	double river_POC02_01(river_time, river) ;
		river_POC02_01:long_name = "river runoff POC02_01" ;
		river_POC02_01:units = "umol L-1" ;
		river_POC02_01:time = "river_time" ;
	double river_POC03_01(river_time, river) ;
		river_POC03_01:long_name = "river runoff POC03_01" ;
		river_POC03_01:units = "umol L-1" ;
		river_POC03_01:time = "river_time" ;
	double river_PON01_01(river_time, river) ;
		river_PON01_01:long_name = "river runoff PON01_01" ;
		river_PON01_01:units = "umol L-1" ;
		river_PON01_01:time = "river_time" ;
	double river_PON02_01(river_time, river) ;
		river_PON02_01:long_name = "river runoff PON02_01" ;
		river_PON02_01:units = "umol L-1" ;
		river_PON02_01:time = "river_time" ;
	double river_PON03_01(river_time, river) ;
		river_PON03_01:long_name = "river runoff PON03_01" ;
		river_PON03_01:units = "umol L-1" ;
		river_PON03_01:time = "river_time" ;
	double river_POP01_01(river_time, river) ;
		river_POP01_01:long_name = "river runoff POP01_01" ;
		river_POP01_01:units = "umol L-1" ;
		river_POP01_01:time = "river_time" ;
	double river_POP02_01(river_time, river) ;
		river_POP02_01:long_name = "river runoff POP02_01" ;
		river_POP02_01:units = "umol L-1" ;
		river_POP02_01:time = "river_time" ;
	double river_POP03_01(river_time, river) ;
		river_POP03_01:long_name = "river runoff POP03_01" ;
		river_POP03_01:units = "umol L-1" ;
		river_POP03_01:time = "river_time" ;

// global attributes:
		:type = "ROMS FORCING file" ;
		:title = "TokyoBay River Forcing" ;
		:grd_file = "TokyoBay2_grid_v3.1.nc" ;
		:rivers = "(1)Edogawa river, (2)Aragawa river (3)Tamagawa river, (4)Nakagawa river,(5)Sumidagawa river, (6)Tsurumigawa river, (7)Obitsugawa river, (8)Yoro river, (9)Koito river" ;
}
